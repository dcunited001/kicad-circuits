.title KiCad schematic
.include "/data/edu/vwcc/etr237/kicad/circuits/spice/KiCad-Spice-Library/Models/Transistor/BJT/BC546.lib"
Cin1 0 Net-_Cin1-Pad2_ 10u
Cout1 out 0 10u
R1 0 Net-_R1-Pad2_ 68k
VCC1 Net-_R1-Pad2_ 0 5
Vin1 Net-_Cin1-Pad2_ 0 sin(0 1m 500)
R3 Net-_R1-Pad2_ 0 10k
R2 0 0 10k
RLoad1 0 out 100k
Q1 NC_01 NC_02 NC_03 BC546B
.ac dec 10 10 100k 
.end
